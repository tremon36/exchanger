package include_local_constants;

`define ALPHA_SELECT_HDR 1'b1
`define ALPHA_SELECT_HSNR 1'b0

`define OP_MODE_FIFTH_ORDER 1'b0
`define OP_MODE_DDR 1'b1

endpackage
